* D:\esim\half_sub\half_sub.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 02/04/22 00:11:04

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  Net-_M1-Pad1_ /vin_A /vdd /vdd mosfet_p		
M9  Net-_M1-Pad1_ /vin_A GND GND mosfet_n		
M2  Net-_M2-Pad1_ /vin_A /vdd /vdd mosfet_p		
M3  Net-_M2-Pad1_ /vin_B /vdd /vdd mosfet_p		
M4  /Diff Net-_M1-Pad1_ Net-_M2-Pad1_ /vdd mosfet_p		
M10  /Diff /vin_A Net-_M10-Pad3_ GND mosfet_n		
M12  Net-_M10-Pad3_ /vin_B GND GND mosfet_n		
M11  /Diff Net-_M1-Pad1_ Net-_M11-Pad3_ GND mosfet_n		
M13  Net-_M11-Pad3_ Net-_M13-Pad2_ GND GND mosfet_n		
M6  Net-_M6-Pad1_ /vin_A /vdd /vdd mosfet_p		
M7  /Borrow Net-_M13-Pad2_ Net-_M6-Pad1_ /vdd mosfet_p		
M14  /Borrow /vin_A GND GND mosfet_n		
M15  /Borrow Net-_M13-Pad2_ GND GND mosfet_n		
M8  Net-_M13-Pad2_ /vin_B /vdd /vdd mosfet_p		
M16  Net-_M13-Pad2_ /vin_B GND GND mosfet_n		
M5  /Diff Net-_M13-Pad2_ Net-_M2-Pad1_ /vdd mosfet_p		
U3  /vin_B PORT		
U2  /vin_A PORT		
U4  /Diff PORT		
U5  /Borrow PORT		
U1  /vdd PORT		

.end
